../../sim/hvl/magic_dual_port.sv