VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER contactResistance REAL ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.0025 ;
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER poly
  TYPE MASTERSLICE ;
END poly

LAYER contact
  TYPE CUT ;
  SPACING 0.075 ;
  PROPERTY contactResistance 10.5 ;
END contact

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 0.19 ;
  WIDTH 0.065 ;
  SPACING 0.065 ;

END metal1

LAYER via1
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.065 ;
  PROPERTY contactResistance 5.69 ;
END via1

LAYER metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.19 0.19 ;
  WIDTH 0.07 ;
  SPACING 0.075 ;
  SPACING 0.07 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal2

LAYER via2
  TYPE CUT ;
  SPACING 0.085 ;
  WIDTH 0.07 ;
  PROPERTY contactResistance 11.39 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 0.19 ;
  WIDTH 0.07 ;
  SPACING 0.07 ;
  SPACING 0.07 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal3

LAYER via3
  TYPE CUT ;
  SPACING 0.085 ;
  WIDTH 0.07 ;
  PROPERTY contactResistance 16.73 ;
END via3

LAYER metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.285 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  SPACING 0.14 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal4

LAYER via4
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  PROPERTY contactResistance 21.44 ;
END via4

LAYER metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.285 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  SPACING 0.14 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal5

LAYER via5
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  PROPERTY contactResistance 24.08 ;
END via5

LAYER metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.285 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  SPACING 0.14 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal6

LAYER via6
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  PROPERTY contactResistance 11.39 ;
END via6

LAYER metal7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.855 0.855 ;
  WIDTH 0.4 ;
  SPACING 0.44 ;
  SPACING 0.44 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal7

LAYER via7
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  PROPERTY contactResistance 5.69 ;
END via7

LAYER metal8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.855 0.855 ;
  WIDTH 0.4 ;
  SPACING 0.44 ;
  SPACING 0.44 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal8

LAYER via8
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  PROPERTY contactResistance 16.73 ;
END via8

LAYER metal9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.71 1.71 ;
  WIDTH 0.8 ;
  SPACING 0.8 ;
  SPACING 0.8 SAMENET ;
  RESISTANCE RPERSQ 0.21 ;
END metal9

LAYER via9
  TYPE CUT ;
  SPACING 0.88 ;
  WIDTH 0.8 ;
  PROPERTY contactResistance 21.44 ;
END via9

LAYER metal10
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.71 1.71 ;
  WIDTH 0.4 ;
  SPACING 0.8 ;
  SPACING 0.8 SAMENET ;
  RESISTANCE RPERSQ 0.21 ;
END metal10

VIARULE M2_M1 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END M2_M1

VIARULE M3_M2 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END M3_M2

VIARULE M4_M3 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END M4_M3

VIARULE M5_M4 GENERATE
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M5_M4

VIARULE M6_M5 GENERATE
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M6_M5

VIARULE M7_M6 GENERATE
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER metal7 ;
    ENCLOSURE 0.13 0.13 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M7_M6

VIARULE M8_M7 GENERATE
  LAYER metal7 ;
    ENCLOSURE 0 0 ;
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 0.8 ;
END M8_M7

VIARULE M9_M8 GENERATE
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER metal9 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 0.8 ;
END M9_M8

VIARULE M10_M9 GENERATE
  LAYER metal9 ;
    ENCLOSURE 0 0 ;
  LAYER metal10 ;
    ENCLOSURE 0 0 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.6 BY 1.6 ;
END M10_M9

VIARULE M1_POLY GENERATE
  LAYER poly ;
    ENCLOSURE 0 0 ;
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER contact ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END M1_POLY

VIA M2_M1_via DEFAULT
  LAYER metal1 ;
    RECT -0.0675 -0.0325 0.0675 0.0325 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.035 -0.0675 0.035 0.0675 ;
END M2_M1_via

VIA M3_M2_via DEFAULT
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END M3_M2_via

VIA M4_M3_via DEFAULT
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M4_M3_via

VIA M5_M4_via DEFAULT
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M5_M4_via

VIA M6_M5_via DEFAULT
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M6_M5_via

VIA M7_M6_via DEFAULT
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M7_M6_via

VIA M8_M7_via DEFAULT
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M8_M7_via

VIA M9_M8_via DEFAULT
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END M9_M8_via

VIA M10_M9_via DEFAULT
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER metal10 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END M10_M9_via

VIA M2_M1_viaB DEFAULT
  LAYER metal1 ;
    RECT -0.0675 -0.0325 0.0675 0.0325 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.0675 -0.035 0.0675 0.035 ;
END M2_M1_viaB

VIA M2_M1_viaC DEFAULT
  LAYER metal1 ;
    RECT -0.0325 -0.0675 0.0325 0.0675 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.035 -0.0675 0.035 0.0675 ;
END M2_M1_viaC

VIA M3_M2_viaB DEFAULT
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END M3_M2_viaB

VIA M3_M2_viaC DEFAULT
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END M3_M2_viaC

VIA M4_M3_viaB DEFAULT
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M4_M3_viaB

SITE CoreSite
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.005 BY 1.005 ;
END CoreSite

MACRO and2
  CLASS CORE ;
  ORIGIN -0.325 0.08 ;
  FOREIGN and2 0.325 -0.08 ;
  SIZE 0.875 BY 1.41 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.6575 0.5125 0.7925 0.5825 ;
      LAYER metal1 ;
        RECT 0.6575 0.515 0.7925 0.5825 ;
      LAYER via1 ;
        RECT 0.6925 0.515 0.7575 0.58 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.865 0.51 1 0.58 ;
      LAYER metal1 ;
        RECT 0.865 0.5125 1 0.58 ;
      LAYER via1 ;
        RECT 0.9 0.5125 0.965 0.5775 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.4225 0.62 0.4925 0.755 ;
      LAYER metal1 ;
        RECT 0.4225 0.62 0.49 0.755 ;
        RECT 0.4225 0.265 0.4875 1.165 ;
      LAYER via1 ;
        RECT 0.425 0.655 0.49 0.72 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.325 1.23 1.2 1.43 ;
        RECT 1.055 1.0025 1.12 1.43 ;
        RECT 0.6525 1.0025 0.7175 1.43 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.325 -0.18 1.2 0.02 ;
        RECT 0.6475 -0.18 0.7125 0.43 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.855 0.6975 0.92 1.1625 ;
      RECT 0.555 0.6975 1.135 0.7625 ;
      RECT 1.07 0.2775 1.135 0.7625 ;
      RECT 1.0575 0.265 1.1225 0.475 ;
  END
END and2

MACRO aoi21
  CLASS CORE ;
  ORIGIN 0 0.08 ;
  FOREIGN aoi21 0 -0.08 ;
  SIZE 0.85 BY 1.41 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.06 0.62 0.195 0.69 ;
      LAYER metal1 ;
        RECT 0.06 0.6225 0.1975 0.6875 ;
      LAYER via1 ;
        RECT 0.095 0.6225 0.16 0.6875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.265 0.62 0.4 0.69 ;
      LAYER metal1 ;
        RECT 0.265 0.62 0.4 0.6875 ;
      LAYER via1 ;
        RECT 0.3 0.6225 0.365 0.6875 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.475 0.62 0.61 0.69 ;
      LAYER metal1 ;
        RECT 0.4775 0.62 0.6125 0.685 ;
        RECT 0.475 0.6225 0.61 0.6875 ;
      LAYER via1 ;
        RECT 0.51 0.6225 0.575 0.6875 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.68 0.5825 0.75 0.7175 ;
      LAYER metal1 ;
        RECT 0.6825 0.265 0.7475 1.1625 ;
        RECT 0.0625 0.4425 0.7475 0.5075 ;
        RECT 0.0625 0.265 0.1275 0.5075 ;
      LAYER via1 ;
        RECT 0.6825 0.6175 0.7475 0.6825 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0 1.23 0.85 1.43 ;
        RECT 0.255 1.0025 0.32 1.43 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.18 0.85 0.02 ;
        RECT 0.4575 -0.18 0.5225 0.375 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.0675 0.8625 0.1325 1.165 ;
      RECT 0.4425 0.8625 0.5075 1.1625 ;
      RECT 0.0675 0.8625 0.5075 0.9275 ;
  END
END aoi21

MACRO buf
  CLASS CORE ;
  ORIGIN -0.2775 0.08 ;
  FOREIGN buf 0.2775 -0.08 ;
  SIZE 0.815 BY 1.41 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.7075 0.55 0.8425 0.62 ;
      LAYER metal1 ;
        RECT 0.7075 0.5525 0.8425 0.6175 ;
      LAYER via1 ;
        RECT 0.7425 0.5525 0.8075 0.6175 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.395 0.605 0.465 0.74 ;
      LAYER metal1 ;
        RECT 0.3975 0.265 0.4625 1.165 ;
      LAYER via1 ;
        RECT 0.3975 0.64 0.4625 0.705 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.2775 1.23 1.0925 1.43 ;
        RECT 0.6775 1.0025 0.7425 1.43 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.2825 -0.18 1.0925 0.02 ;
        RECT 0.6725 -0.18 0.7375 0.4025 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.9375 0.265 1.0025 1.165 ;
      RECT 0.56 0.72 1.0025 0.785 ;
  END
END buf

MACRO dff
  CLASS CORE ;
  ORIGIN -0.2225 -0.1125 ;
  FOREIGN dff 0.2225 0.1125 ;
  SIZE 3.89 BY 1.41 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.675 0.7925 0.81 0.8625 ;
      LAYER metal1 ;
        RECT 0.675 0.795 0.81 0.86 ;
      LAYER via1 ;
        RECT 0.71 0.795 0.775 0.86 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 1.14 0.7725 1.275 0.8425 ;
      LAYER metal1 ;
        RECT 1.14 0.775 1.275 0.84 ;
        RECT 1.14 0.4575 1.205 1.355 ;
      LAYER via1 ;
        RECT 1.175 0.775 1.24 0.84 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.9025 0.45 3.9675 1.35 ;
        RECT 3.54 0.94 3.9675 1.005 ;
    END
  END Q
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.2225 1.4225 4.1125 1.6225 ;
        RECT 3.6425 1.1875 3.7075 1.6225 ;
        RECT 2.24 1.195 2.305 1.6225 ;
        RECT 0.6625 1.195 0.7275 1.6225 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.2225 0.0125 4.1125 0.2125 ;
        RECT 3.6375 0.0125 3.7025 0.635 ;
        RECT 2.235 0.0125 2.3 0.5925 ;
        RECT 0.6575 0.0125 0.7225 0.6575 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 2.9525 0.45 3.0175 1.3475 ;
      RECT 2.9525 0.76 3.0875 0.825 ;
      RECT 2.5575 0.4575 2.6225 1.3575 ;
      RECT 2.1375 0.9475 2.6225 1.0125 ;
      RECT 2.3425 0.765 2.4775 0.83 ;
      RECT 2.34 0.7625 2.475 0.8275 ;
      RECT 1.5325 0.4575 1.5975 1.355 ;
      RECT 1.5325 0.7625 1.6675 0.8275 ;
      RECT 0.95 0.3275 1.015 1.3575 ;
      RECT 0.915 1.2175 1.05 1.2825 ;
      RECT 0.915 0.6225 1.05 0.6875 ;
      RECT 3.7 0.76 3.8375 0.825 ;
      RECT 3.3525 0.45 3.4175 1.35 ;
      RECT 3.1375 1.0525 3.2725 1.1175 ;
      RECT 3.1275 0.62 3.2625 0.685 ;
      RECT 2.72 0.6225 2.855 0.6875 ;
      RECT 2.7 1.06 2.835 1.125 ;
      RECT 1.9575 0.4575 2.0225 1.3575 ;
      RECT 1.725 1.06 1.86 1.125 ;
      RECT 1.7075 0.6225 1.8425 0.6875 ;
      RECT 1.2925 0.6225 1.4275 0.6875 ;
      RECT 1.2725 0.9675 1.4075 1.0325 ;
      RECT 0.4525 0.6225 0.5875 0.6875 ;
      RECT 0.29 0.37 0.355 1.3575 ;
    LAYER metal2 ;
      RECT 3.1375 1.05 3.2725 1.12 ;
      RECT 3.145 0.8975 3.215 1.12 ;
      RECT 2.785 0.8975 3.215 0.9675 ;
      RECT 2.785 0.62 2.855 0.9675 ;
      RECT 1.7075 0.62 2.855 0.69 ;
      RECT 1.74 0.37 1.81 0.69 ;
      RECT 0.2875 0.37 0.3575 0.505 ;
      RECT 0.2875 0.37 1.81 0.44 ;
      RECT 0.915 1.215 1.81 1.285 ;
      RECT 1.74 1.0575 1.81 1.285 ;
      RECT 1.725 1.0575 2.835 1.1275 ;
      RECT 0.2875 0.965 1.4075 1.035 ;
      RECT 0.2875 0.9 0.3575 1.035 ;
      RECT 2.9525 0.7575 3.835 0.8275 ;
      RECT 3.1275 0.6175 3.2625 0.6875 ;
      RECT 1.5325 0.76 2.475 0.83 ;
      RECT 0.4525 0.62 1.4275 0.69 ;
    LAYER via1 ;
      RECT 3.735 0.76 3.8 0.825 ;
      RECT 3.1725 1.0525 3.2375 1.1175 ;
      RECT 3.1625 0.62 3.2275 0.685 ;
      RECT 2.9875 0.76 3.0525 0.825 ;
      RECT 2.755 0.6225 2.82 0.6875 ;
      RECT 2.735 1.06 2.8 1.125 ;
      RECT 2.375 0.7625 2.44 0.8275 ;
      RECT 1.76 1.06 1.825 1.125 ;
      RECT 1.7425 0.6225 1.8075 0.6875 ;
      RECT 1.5675 0.7625 1.6325 0.8275 ;
      RECT 1.3275 0.6225 1.3925 0.6875 ;
      RECT 1.3075 0.9675 1.3725 1.0325 ;
      RECT 0.95 0.6225 1.015 0.6875 ;
      RECT 0.95 1.2175 1.015 1.2825 ;
      RECT 0.4875 0.6225 0.5525 0.6875 ;
      RECT 0.29 0.405 0.355 0.47 ;
      RECT 0.29 0.935 0.355 1 ;
  END
END dff

MACRO inv
  CLASS CORE ;
  ORIGIN -0.0675 0.08 ;
  FOREIGN inv 0.0675 -0.08 ;
  SIZE 0.41 BY 1.4075 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.13 0.55 0.265 0.62 ;
      LAYER metal1 ;
        RECT 0.13 0.5525 0.265 0.6175 ;
      LAYER via1 ;
        RECT 0.165 0.5525 0.23 0.6175 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.3375 0.605 0.4075 0.74 ;
      LAYER metal1 ;
        RECT 0.3375 0.605 0.405 0.74 ;
        RECT 0.3375 0.265 0.4025 1.165 ;
      LAYER via1 ;
        RECT 0.34 0.64 0.405 0.705 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.0675 1.23 0.4775 1.43 ;
        RECT 0.135 1.0025 0.2 1.43 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.0675 -0.18 0.4775 0.02 ;
        RECT 0.13 -0.18 0.195 0.4025 ;
    END
  END vss!
END inv

MACRO latch
  CLASS CORE ;
  ORIGIN -0.35 -0.105 ;
  FOREIGN latch 0.35 0.105 ;
  SIZE 2.44 BY 1.41 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 1.265 0.765 1.4 0.835 ;
      LAYER metal1 ;
        RECT 1.265 0.7675 1.4 0.8325 ;
        RECT 1.265 0.45 1.33 1.3475 ;
      LAYER via1 ;
        RECT 1.3 0.7675 1.365 0.8325 ;
    END
  END D
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.83 0.73 0.965 0.795 ;
    END
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 1.6575 0.795 2.5025 0.865 ;
      LAYER metal1 ;
        RECT 2.37 0.8 2.505 0.865 ;
        RECT 2.3675 0.7975 2.5025 0.8625 ;
        RECT 1.6575 0.7975 1.7925 0.8625 ;
        RECT 1.6575 0.45 1.7225 1.3475 ;
      LAYER via1 ;
        RECT 1.6925 0.7975 1.7575 0.8625 ;
        RECT 2.4025 0.7975 2.4675 0.8625 ;
    END
  END Q
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.35 1.415 2.79 1.615 ;
        RECT 2.3225 1.1875 2.3875 1.615 ;
        RECT 0.7575 1.1875 0.8225 1.615 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.35 0.005 2.79 0.205 ;
        RECT 2.3175 0.005 2.3825 0.585 ;
        RECT 0.7525 0.005 0.8175 0.5925 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 2.5925 0.45 2.6575 1.35 ;
      RECT 2.22 0.94 2.6575 1.005 ;
      RECT 1.0875 0.32 1.1525 1.35 ;
      RECT 1.0625 0.325 1.1975 0.39 ;
      RECT 0.4175 0.37 0.4825 1.35 ;
      RECT 0.4175 0.615 0.555 0.68 ;
      RECT 2.0475 0.45 2.1125 1.35 ;
      RECT 1.825 1.0525 1.96 1.1175 ;
      RECT 1.815 0.62 1.95 0.685 ;
      RECT 1.4175 0.615 1.5525 0.68 ;
      RECT 1.3975 1.0525 1.5325 1.1175 ;
      RECT 0.595 1.0525 0.73 1.1175 ;
    LAYER metal2 ;
      RECT 0.42 1.22 1.895 1.29 ;
      RECT 1.825 1.05 1.895 1.29 ;
      RECT 0.42 0.6125 0.49 1.29 ;
      RECT 1.825 1.05 1.96 1.12 ;
      RECT 0.42 0.6125 1.5525 0.6825 ;
      RECT 1.815 0.6175 1.95 0.6875 ;
      RECT 1.8325 0.3225 1.9025 0.6875 ;
      RECT 1.0625 0.3225 1.9025 0.3925 ;
      RECT 0.595 1.05 1.5325 1.12 ;
      RECT 1.085 0.985 1.155 1.12 ;
    LAYER via1 ;
      RECT 1.86 1.0525 1.925 1.1175 ;
      RECT 1.85 0.62 1.915 0.685 ;
      RECT 1.4525 0.615 1.5175 0.68 ;
      RECT 1.4325 1.0525 1.4975 1.1175 ;
      RECT 1.0975 0.325 1.1625 0.39 ;
      RECT 1.0875 1.02 1.1525 1.085 ;
      RECT 0.63 1.0525 0.695 1.1175 ;
      RECT 0.455 0.615 0.52 0.68 ;
  END
END latch

MACRO mux2
  CLASS CORE ;
  ORIGIN 0.385 0.08 ;
  FOREIGN mux2 -0.385 -0.08 ;
  SIZE 2.0325 BY 1.41 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.66 0.54 0.795 0.61 ;
      LAYER metal1 ;
        RECT 0.66 0.54 0.795 0.6075 ;
      LAYER via1 ;
        RECT 0.695 0.5425 0.76 0.6075 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 1.28 0.68 1.415 0.75 ;
      LAYER metal1 ;
        RECT 1.28 0.6825 1.415 0.7475 ;
        RECT 1.2775 0.685 1.4125 0.75 ;
      LAYER via1 ;
        RECT 1.315 0.6825 1.38 0.7475 ;
    END
  END B
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.17 0.6825 1.21 0.7525 ;
      LAYER metal1 ;
        RECT 1.075 0.685 1.21 0.75 ;
        RECT 0.17 0.685 0.305 0.75 ;
      LAYER via1 ;
        RECT 0.205 0.685 0.27 0.75 ;
        RECT 1.11 0.685 1.175 0.75 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT -0.2975 0.605 -0.2275 0.74 ;
      LAYER metal1 ;
        RECT -0.295 0.265 -0.23 1.165 ;
      LAYER via1 ;
        RECT -0.295 0.64 -0.23 0.705 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.385 1.23 1.6475 1.43 ;
        RECT 0.8525 1.0025 0.9175 1.43 ;
        RECT 0.0725 1.0025 0.1375 1.43 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT -0.385 -0.18 1.6475 0.02 ;
        RECT 1.055 -0.18 1.12 0.36 ;
        RECT 0.0625 -0.18 0.1275 0.4025 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 1.275 0.815 1.34 1.0325 ;
      RECT 1.275 0.815 1.5475 0.88 ;
      RECT 1.4825 0.2675 1.5475 0.88 ;
      RECT 1.4125 0.2675 1.5475 0.3325 ;
      RECT 0.665 0.8625 0.73 1.165 ;
      RECT 1.04 1.0975 1.54 1.1625 ;
      RECT 1.475 0.9475 1.54 1.1625 ;
      RECT 1.04 0.8625 1.105 1.1625 ;
      RECT 0.665 0.8625 1.105 0.9275 ;
      RECT 0.425 0.265 0.49 1.165 ;
      RECT 0.425 0.685 0.995 0.75 ;
      RECT 0.66 0.265 0.725 0.425 ;
      RECT 0.66 0.2675 0.795 0.3325 ;
      RECT -0.0925 0.625 0.0425 0.69 ;
    LAYER metal2 ;
      RECT -0.0925 0.6225 0.0425 0.6925 ;
      RECT -0.055 0.265 0.015 0.6925 ;
      RECT -0.0575 0.265 1.5475 0.335 ;
    LAYER via1 ;
      RECT 1.4475 0.2675 1.5125 0.3325 ;
      RECT 0.695 0.2675 0.76 0.3325 ;
      RECT -0.0575 0.625 0.0075 0.69 ;
  END
END mux2

MACRO nand2
  CLASS CORE ;
  ORIGIN 0 0.08 ;
  FOREIGN nand2 0 -0.08 ;
  SIZE 0.6 BY 1.41 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.0725 0.5125 0.2075 0.5825 ;
      LAYER metal1 ;
        RECT 0.0725 0.515 0.2075 0.5825 ;
      LAYER via1 ;
        RECT 0.1075 0.515 0.1725 0.58 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.28 0.51 0.415 0.58 ;
      LAYER metal1 ;
        RECT 0.28 0.5125 0.415 0.58 ;
      LAYER via1 ;
        RECT 0.315 0.5125 0.38 0.5775 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.2675 0.805 0.3375 0.94 ;
      LAYER metal1 ;
        RECT 0.27 0.65 0.555 0.715 ;
        RECT 0.49 0.2775 0.555 0.715 ;
        RECT 0.4725 0.265 0.5375 0.475 ;
        RECT 0.27 0.65 0.335 1.165 ;
      LAYER via1 ;
        RECT 0.27 0.84 0.335 0.905 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0 1.23 0.6 1.43 ;
        RECT 0.47 1.0025 0.535 1.43 ;
        RECT 0.0675 1.0025 0.1325 1.43 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.18 0.6 0.02 ;
        RECT 0.0625 -0.18 0.1275 0.43 ;
    END
  END vss!
END nand2

MACRO nor2
  CLASS CORE ;
  ORIGIN 0 0.08 ;
  FOREIGN nor2 0 -0.08 ;
  SIZE 0.6 BY 1.41 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.0725 0.645 0.2075 0.715 ;
      LAYER metal1 ;
        RECT 0.0725 0.6475 0.2075 0.7125 ;
      LAYER via1 ;
        RECT 0.1075 0.6475 0.1725 0.7125 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.28 0.6425 0.415 0.7125 ;
      LAYER metal1 ;
        RECT 0.28 0.645 0.415 0.7125 ;
      LAYER via1 ;
        RECT 0.315 0.645 0.38 0.71 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.4275 0.4875 0.5625 0.5575 ;
      LAYER metal1 ;
        RECT 0.4975 0.49 0.5625 1.065 ;
        RECT 0.47 0.8975 0.535 1.165 ;
        RECT 0.2725 0.4925 0.5625 0.5575 ;
        RECT 0.4275 0.49 0.5625 0.5575 ;
        RECT 0.2725 0.265 0.3375 0.5575 ;
      LAYER via1 ;
        RECT 0.4625 0.49 0.5275 0.555 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0 1.23 0.6 1.43 ;
        RECT 0.0675 1.0025 0.1325 1.43 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.18 0.6 0.02 ;
        RECT 0.475 -0.18 0.54 0.4025 ;
        RECT 0.0625 -0.18 0.1275 0.4 ;
    END
  END vss!
END nor2

MACRO oai21
  CLASS CORE ;
  ORIGIN 0 0.08 ;
  FOREIGN oai21 0 -0.08 ;
  SIZE 0.82 BY 1.41 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.065 0.595 0.2 0.665 ;
      LAYER metal1 ;
        RECT 0.0625 0.5975 0.2 0.6625 ;
      LAYER via1 ;
        RECT 0.1 0.5975 0.165 0.6625 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.27 0.5975 0.405 0.6675 ;
      LAYER metal1 ;
        RECT 0.27 0.6 0.405 0.665 ;
      LAYER via1 ;
        RECT 0.305 0.6 0.37 0.665 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.4775 0.5975 0.6125 0.6675 ;
      LAYER metal1 ;
        RECT 0.4775 0.6 0.6125 0.665 ;
      LAYER via1 ;
        RECT 0.5125 0.6 0.5775 0.665 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.4425 0.7825 0.5775 0.8525 ;
      LAYER metal1 ;
        RECT 0.4425 0.785 0.7475 0.85 ;
        RECT 0.6825 0.265 0.7475 0.85 ;
        RECT 0.4425 0.785 0.5075 1.1325 ;
      LAYER via1 ;
        RECT 0.4775 0.785 0.5425 0.85 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0 1.23 0.82 1.43 ;
        RECT 0.6825 0.99 0.7475 1.43 ;
        RECT 0.0675 0.9875 0.1325 1.43 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.18 0.82 0.02 ;
        RECT 0.255 -0.18 0.32 0.375 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.0625 0.44 0.5225 0.505 ;
      RECT 0.4575 0.265 0.5225 0.505 ;
      RECT 0.0625 0.265 0.1275 0.505 ;
  END
END oai21

MACRO or2
  CLASS CORE ;
  ORIGIN -0.3225 0.08 ;
  FOREIGN or2 0.3225 -0.08 ;
  SIZE 0.8525 BY 1.41 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.6375 0.69 0.7725 0.76 ;
      LAYER metal1 ;
        RECT 0.6375 0.6925 0.7725 0.7575 ;
      LAYER via1 ;
        RECT 0.6725 0.6925 0.7375 0.7575 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.845 0.69 0.98 0.76 ;
      LAYER metal1 ;
        RECT 0.845 0.6925 0.98 0.7575 ;
      LAYER via1 ;
        RECT 0.88 0.6925 0.945 0.7575 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.385 0.6 0.455 0.735 ;
      LAYER metal1 ;
        RECT 0.3875 0.265 0.4525 1.165 ;
      LAYER via1 ;
        RECT 0.3875 0.635 0.4525 0.7 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.3225 1.23 1.17 1.43 ;
        RECT 0.6325 1.0025 0.6975 1.43 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.3225 -0.18 1.175 0.02 ;
        RECT 1.0375 -0.18 1.1025 0.4025 ;
        RECT 0.6275 -0.18 0.6925 0.3975 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 1.035 0.94 1.1 1.165 ;
      RECT 1.055 0.4925 1.12 1.14 ;
      RECT 0.525 0.4925 1.12 0.5575 ;
      RECT 0.835 0.265 0.9 0.5575 ;
  END
END or2

MACRO xnor2
  CLASS CORE ;
  ORIGIN -0.0725 -0.1 ;
  FOREIGN xnor2 0.0725 0.1 ;
  SIZE 1.395 BY 1.41 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.1425 0.8725 1.175 0.9425 ;
      LAYER metal1 ;
        RECT 1.04 0.875 1.175 0.94 ;
        RECT 0.1425 0.875 0.2775 0.94 ;
      LAYER via1 ;
        RECT 0.1775 0.875 0.2425 0.94 ;
        RECT 1.075 0.875 1.14 0.94 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.48 0.7325 0.9625 0.8025 ;
      LAYER metal1 ;
        RECT 0.8275 0.735 0.9625 0.8 ;
        RECT 0.48 0.735 0.615 0.8 ;
        RECT 0.4775 0.7325 0.6125 0.7975 ;
      LAYER via1 ;
        RECT 0.515 0.735 0.58 0.8 ;
        RECT 0.8625 0.735 0.9275 0.8 ;
    END
  END B
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.0725 1.41 1.4675 1.61 ;
        RECT 1.2475 1.0925 1.3125 1.61 ;
        RECT 0.5425 1.145 0.6075 1.61 ;
        RECT 0.14 1.1825 0.205 1.61 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.0725 0 1.4675 0.2 ;
        RECT 0.5475 0 0.6125 0.4875 ;
    END
  END vss!
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.82 1.1325 1.3975 1.2025 ;
        RECT 1.3275 0.5525 1.3975 1.2025 ;
        RECT 1.035 0.5525 1.3975 0.6225 ;
        RECT 1.035 0.265 1.105 0.6225 ;
        RECT 0.82 1.1325 0.89 1.2675 ;
      LAYER metal1 ;
        RECT 1.0375 0.265 1.1025 0.4025 ;
        RECT 0.8225 1.125 0.8875 1.3075 ;
      LAYER via1 ;
        RECT 0.8225 1.1675 0.8875 1.2325 ;
        RECT 1.0375 0.3 1.1025 0.365 ;
    END
  END Y
  OBS
    LAYER metal1 ;
      RECT 0.8225 0.4675 1.3125 0.5325 ;
      RECT 1.2475 0.31 1.3125 0.5325 ;
      RECT 0.8225 0.315 0.8875 0.5325 ;
      RECT 0.3475 0.5875 0.4125 1.3425 ;
      RECT 0.135 0.5875 0.7625 0.6525 ;
      RECT 0.135 0.285 0.2 0.6525 ;
  END
END xnor2

MACRO xor2
  CLASS CORE ;
  ORIGIN -0.0825 0.08 ;
  FOREIGN xor2 0.0825 -0.08 ;
  SIZE 1.42 BY 1.41 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.1525 0.6925 1.2 0.7625 ;
      LAYER metal1 ;
        RECT 1.065 0.695 1.21 0.76 ;
        RECT 0.1525 0.695 0.2875 0.76 ;
      LAYER via1 ;
        RECT 0.1875 0.695 0.2525 0.76 ;
        RECT 1.1 0.695 1.165 0.76 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.4875 0.5475 1.0075 0.6175 ;
      LAYER metal1 ;
        RECT 0.8725 0.55 1.0075 0.615 ;
        RECT 0.4875 0.55 0.6225 0.615 ;
      LAYER via1 ;
        RECT 0.5225 0.55 0.5875 0.615 ;
        RECT 0.9075 0.55 0.9725 0.615 ;
    END
  END B
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.0825 1.23 1.5025 1.43 ;
        RECT 0.5525 1.0025 0.6175 1.43 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.0825 -0.18 1.5025 0.02 ;
        RECT 1.2825 -0.18 1.3475 0.295 ;
        RECT 0.5575 -0.18 0.6225 0.2675 ;
        RECT 0.145 -0.18 0.21 0.265 ;
    END
  END vss!
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 1.055 0.9775 1.35 1.0475 ;
        RECT 1.28 0.3225 1.35 1.0475 ;
        RECT 0.855 0.3225 1.35 0.3925 ;
        RECT 1.055 0.975 1.125 1.11 ;
        RECT 0.855 0.135 0.925 0.3925 ;
      LAYER metal1 ;
        RECT 1.0575 0.975 1.1225 1.165 ;
        RECT 0.8575 0.13 0.9225 0.2725 ;
      LAYER via1 ;
        RECT 0.8575 0.17 0.9225 0.235 ;
        RECT 1.0575 1.01 1.1225 1.075 ;
    END
  END Y
  OBS
    LAYER metal1 ;
      RECT 1.2825 0.8375 1.3475 1.1625 ;
      RECT 0.855 0.8375 0.92 1.1525 ;
      RECT 0.855 0.8375 1.3475 0.9025 ;
      RECT 0.1525 0.85 0.2175 1.165 ;
      RECT 0.1525 0.85 0.4175 0.915 ;
      RECT 0.3525 0.13 0.4175 0.915 ;
      RECT 0.3525 0.4125 0.8 0.4775 ;
  END
END xor2

END LIBRARY
